`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:31:51 10/22/2018 
// Design Name: 
// Module Name:    Combinacional4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module Combinacional4(
    input [2:0]Q,
    output [2:0]Qnext
    );

	assign Qnext = Q+1;
	
						
endmodule
