`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:41:12 09/24/2018 
// Design Name: 
// Module Name:    Decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Decoder(
    input [3:0] A,
    output [6:0] Seg
    );

	assign Seg =	(A==4'b0000)? 7'b1000000://0
						(A==4'b0001)? 7'b1111001://1
						(A==4'b0010)? 7'b0100100://2
						(A==4'b0011)? 7'b0110000://3
						(A==4'b0100)? 7'b0011001://4
						(A==4'b0101)? 7'b0010010://5
						(A==4'b0110)? 7'b0000010://6
						(A==4'b0111)? 7'b1111000://7
						(A==4'b1000)? 7'b0000000://8
						(A==4'b1001)? 7'b0011000://9
						(A==4'b1010)? 7'b0001000://A
						(A==4'b1011)? 7'b0000011://B
						(A==4'b1100)? 7'b1000110://C
						(A==4'b1101)? 7'b0100001://D
						(A==4'b1110)? 7'b0000110://E
						(A==4'b1111)? 7'b0001110://F
													  0;

endmodule
